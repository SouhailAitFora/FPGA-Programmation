module test_MED;

logic BYP,DSI,CLK ;
logic [7:0] DI,DO ;
logic [7:0] LIST_TEST [8:0] ;
logic [7:0] LIST_TEST [8:0] ;



 

MED MED1(.BYP(BYP)  ,.DSI(DSI),  .CLK(CLK),  .DI(DI),  .DO(DO));













endmodule